
localparam adder_unsigned     = 2'b00;
localparam adder_1sComplement = 2'b01;
localparam adder_2sComplement = 2'b10;
